module tics_module_name(out_2, out_6, in_5, in_4, in_7, in_3);
  output out_2;
  output out_6;
  input in_3;
  input in_4;
  input in_5;
  input in_7;
  supply0 gnd;
  wire wire_8;
  wire wire_9;
  wire wire_10;
  wire wire_11;
  pullup plu_2(out_2);
  pullup plu_6(out_6);
  pullup plu_9(wire_9);
  pullup plu_8(wire_8);
  pullup plu_11(wire_11);
  pullup plu_10(wire_10);
  pullup plu_2(out_2);
  pullup plu_6(out_6);
  nmos mos_1(out_2, gnd, out_6);
  nmos mos_2(out_6, gnd, wire_8);
  nmos mos_3(out_6, gnd, in_5);
  nmos mos_4(wire_9, gnd, in_5);
  nmos mos_5(wire_9, gnd, wire_8);
  nmos mos_6(wire_8, gnd, wire_9);
  nmos mos_7(wire_9, gnd, wire_10);
  nmos mos_8(out_6, gnd, out_2);
  nmos mos_9(wire_8, gnd, in_4);
  nmos mos_10(wire_8, gnd, in_3);
  nmos mos_11(wire_11, gnd, in_4);
  nmos mos_12(wire_11, gnd, wire_8);
  nmos mos_13(wire_11, gnd, wire_10);
  nmos mos_14(out_6, gnd, out_2);
  nmos mos_15(out_2, gnd, wire_11);
  nmos mos_16(wire_10, gnd, wire_11);
  nmos mos_17(out_2, gnd, out_6);
  nmos mos_18(wire_10, gnd, in_3);
  nmos mos_19(wire_10, gnd, in_7);
  nmos mos_21(out_2, gnd, in_3);
endmodule
